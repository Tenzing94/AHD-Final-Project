----------------------------------------------------------------------------------
-- Company: NYU Tandon AHD
-- Engineer: 
-- 
-- Create Date: 11/05/2018 02:34:14 PM
-- Design Name: 
-- Module Name: imem - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Revision 0.02 - Tenzing - I changed line 40 from '(31 downto 2)' to '(31 downto 0)'
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

entity imem is
    Port ( 
           in_pc : in std_logic_vector (31 downto 0);
           out_imem : out std_logic_vector (31 downto 0));
end imem;

architecture Behavioral of imem is
    -- ROM: Instruction Memory -- 
    type ROM_type is array (0 to 503) of std_logic_vector(7 downto 0);
     constant rom_data: ROM_type:=(
              "00000000","00000000","00000000","00000011",
     "00000000","00100001","00001000","00000011",
     "00000000","01000010","00010000","00000011",
     "00000000","01100011","00011000","00000011",
     "00000000","10000100","00100000","00000011",
     "00011100","00000011","00000000","00111000",
     "00011100","00000100","00000000","00111000",
     "00010100","01100011","00000000","00001000",
     "00000000","01100100","00011000","00000111",
     "00000000","10000100","00100000","00000011",
     "00011100","00000001","00000000","00110100",
     "00010100","00100001","00000000","00010000",
     "00011100","10000100","00000000","00110101",
     "00000000","10000011","00100000","00000101",
     "00000000","00100100","00001000","00000111",
     "00000000","10000100","00100000","00000011",
     "00011100","00000010","00000000","00110110",
     "00010100","01000010","00000000","00010000",
     "00011100","10000100","00000000","00110111",
     "00000000","10000011","00100000","00000101",
     "00000000","01000100","00010000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","10100101","00101000","00000011",
     "00000100","10100101","00000000","00000100",
     "00011100","00000110","00000000","00000000",
     "00010100","11000110","00000000","00010000",
     "00011100","00000100","00000000","00000001",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","00100110","00001000","00000001",
     "00011100","00000110","00000000","00000010",
     "00010100","11000110","00000000","00010000",
     "00011100","00000100","00000000","00000011",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","01000110","00010000","00000001",
     "00000000","00100010","00001000","00000001",
     "00000000","11100111","00111000","00000011",
     "00000100","11100111","00000000","00001011",
     "00000010","00010000","10000000","00000011",
     "00000010","00110001","10001000","00000011",
     "00000000","00100010","10000000","00000101",
     "00000000","00100010","10001000","00001001",
     "00000010","00010001","00001000","00001001",
     "00000001","01101011","01011000","00000011",
     "00000001","01100010","01011000","00000111",
     "00000001","10001100","01100000","00000011",
     "00000001","10000001","01100000","00000111",
     "00000001","11001110","01110000","00000011",
     "00000001","11001011","01110000","00000111",
     "00000001","11101111","01111000","00000011",
     "00000001","11101100","01111000","00000111",
     "00001101","01101011","00000000","00011111",
     "00001101","11001110","00000000","00011111",
     "00101000","00001110","00000000","00000011",
     "00010101","11101111","00000000","00000001",
     "00001001","11001110","00000000","00000001",
     "00101101","11000000","11111111","11111101",
     "00000001","01001010","01010000","00000011",
     "00101001","01100000","00000000","00000111",
     "00010101","01001010","00000000","00000001",
     "00100101","10000000","00000000","00000011",
     "00010101","10001100","00000000","00000001",
     "00001001","01101011","00000000","00000001",
     "00110000","00000000","00000000","00111101",
     "00010001","01001010","00000000","00000001",
     "00110000","00000000","00000000","01000000",
     "00000001","10001100","01100000","00000011",
     "00000001","10001010","01100000","00000111",
     "00000001","10001111","01100000","00000111",
     "00000000","00100001","00001000","00000011",
     "00000000","00101100","00001000","00000111",
     "00011100","10100110","00000000","00000000",
     "00010100","11000110","00000000","00010000",
     "00000100","10100101","00000000","00000001",
     "00011100","10100100","00000000","00000000",
     "00000100","10100101","00000000","00000001",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","00100110","00001000","00000001",
     "00000010","00010000","10000000","00000011",
     "00000010","00110001","10001000","00000011",
     "00000000","00100010","10000000","00000101",
     "00000000","00100010","10001000","00001001",
     "00000010","00010001","00010000","00001001",
     "00000001","01101011","01011000","00000011",
     "00000001","01100001","01011000","00000111",
     "00000001","10001100","01100000","00000011",
     "00000001","10000010","01100000","00000111",
     "00000001","11001110","01110000","00000011",
     "00000001","11001011","01110000","00000111",
     "00000001","11101111","01111000","00000011",
     "00000001","11101100","01111000","00000111",
     "00001101","01101011","00000000","00011111",
     "00001101","11001110","00000000","00011111",
     "00101000","00001110","00000000","00000011",
     "00010101","11101111","00000000","00000001",
     "00001001","11001110","00000000","00000001",
     "00101101","11000000","11111111","11111101",
     "00000001","01001010","01010000","00000011",
     "00101001","01100000","00000000","00000111",
     "00010101","01001010","00000000","00000001",
     "00100101","10000000","00000000","00000011",
     "00010101","10001100","00000000","00000001",
     "00001001","01101011","00000000","00000001",
     "00110000","00000000","00000000","01100111",
     "00010001","01001010","00000000","00000001",
     "00110000","00000000","00000000","01101010",
     "00000001","10001100","01100000","00000011",
     "00000001","10001010","01100000","00000111",
     "00000001","10001111","01100000","00000111",
     "00000000","01000010","00010000","00000011",
     "00000000","01001100","00010000","00000111",
     "00011100","10100110","00000000","00000000",
     "00010100","11000110","00000000","00010000",
     "00000100","10100101","00000000","00000001",
     "00011100","10100100","00000000","00000000",
     "00000100","10100101","00000000","00000001",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","01000110","00010000","00000001",
     "11111100","00000000","00000000","00000000"
      );  
    begin
        out_imem <= rom_data(to_integer(unsigned(in_pc(31 downto 0)))) & rom_data(to_integer(unsigned(in_pc(31 downto 0)) + 1 )) & rom_data(to_integer(unsigned(in_pc(31 downto 0)) + 2 )) & rom_data(to_integer(unsigned(in_pc(31 downto 0)) + 3 ));
end Behavioral;

