----------------------------------------------------------------------------------
-- Company: NYU Tandon AHD
-- Engineer: 
-- 
-- Create Date: 11/05/2018 02:34:14 PM
-- Design Name: 
-- Module Name: imem - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Revision 0.02 - Tenzing - I changed line 40 from '(31 downto 2)' to '(31 downto 0)'
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

entity imem is
    Port ( 
           in_pc : in std_logic_vector (31 downto 0);
           out_imem : out std_logic_vector (31 downto 0));
end imem;

architecture Behavioral of imem is
    -- ROM: Instruction Memory -- 
    type ROM_type is array (0 to 111) of std_logic_vector(7 downto 0);
     constant rom_data: ROM_type:=(
              "00000000","00000000","00000000","00000011",
     "00000001","01101011","01011000","00000011",
     "00000001","01100010","01011000","00000111",
     "00000001","10001100","01100000","00000011",
     "00000001","10000001","01100000","00000111",
     "00000001","11001110","01110000","00000011",
     "00000001","11001011","01110000","00000111",
     "00000001","11101111","01111000","00000011",
     "00000001","11101100","01111000","00000111",
     "00001101","01101011","00000000","00011111",
     "00001101","11001110","00000000","00011111",
     "00101000","00001110","00000000","00000011",
     "00010101","11101111","00000000","00000001",
     "00001001","11001110","00000000","00000001",
     "00101101","11000000","11111111","11111101",
     "00000001","01001010","01010000","00000011",
     "00101001","01100000","00000000","00000111",
     "00010101","01001010","00000000","00000001",
     "00100101","10000000","00000000","00000011",
     "00010101","10001100","00000000","00000001",
     "00001001","01101011","00000000","00000001",
     "00110000","00000000","00000000","00010000",
     "00010001","01001010","00000000","00000001",
     "00110000","00000000","00000000","00010011",
     "00000001","10001100","01100000","00000011",
     "00000001","10001010","01100000","00000111",
     "00000001","10001111","01100000","00000111",
     "11111100","00000000","00000000","00000000"
      );  
    begin
        out_imem <= rom_data(to_integer(unsigned(in_pc(31 downto 0)))) & rom_data(to_integer(unsigned(in_pc(31 downto 0)) + 1 )) & rom_data(to_integer(unsigned(in_pc(31 downto 0)) + 2 )) & rom_data(to_integer(unsigned(in_pc(31 downto 0)) + 3 ));
end Behavioral;

