----------------------------------------------------------------------------------
-- Company: NYU Tandon AHD
-- Engineer: 
-- 
-- Create Date: 11/06/2018
-- Design Name: 
-- Module Name: rf - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: Register File for MIPS32-AHD 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created (11/06/2018 12:09PM)
-- Revision 0.02 - Corrected some typos. (11/06/2018 12:11PM)
-- Revision 0.03 - Wrote the body of the rf. (11/06/2018 12:50PM)
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

entity rf is
    Port (
            CLK, WE3   : in std_logic;
            A1, A2, A3 : in std_logic_vector(4 downto 0);
            WD3        : in std_logic_vector(31 downto 0);   
            RD1, RD2   : out std_logic_vector(31 downto 0)
    );
end rf;

architecture Behavioral of rf is

type Register_Type is array (0 to 31) of std_logic_vector(31 downto 0);

signal Reg32 : Register_Type := (
    "00000000000000000000000000000000", "10000000000000001000000000000000",
    "00000000000000000000000000000001", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000",
    "00000000000000000000000000000000", "00000000000000000000000000000000"
);

begin

    -- write
    process(CLK)
    begin
        if(rising_edge(CLK) AND WE3 = '1') then
            Reg32(to_integer(unsigned(A3))) <= WD3;
        end if;   
    end process;
    
    -- read
    RD1 <= Reg32(to_integer(unsigned(A1)));
    RD2 <= Reg32(to_integer(unsigned(A2)));
    


end Behavioral;
