----------------------------------------------------------------------------------
-- Company: NYU Tandon AHD
-- Engineer: 
-- 
-- Create Date: 11/05/2018 02:34:14 PM
-- Design Name: 
-- Module Name: imem - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Revision 0.02 - Tenzing - I changed line 40 from '(31 downto 2)' to '(31 downto 0)'
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

entity imem is
    Port ( 
           in_pc : in std_logic_vector (31 downto 0);
           out_imem : out std_logic_vector (31 downto 0));
end imem;

architecture Behavioral of imem is
    -- ROM: Instruction Memory -- 
    type ROM_type is array (0 to 1887) of std_logic_vector(7 downto 0);
     constant rom_data: ROM_type:=(
            "00000000","01100011","00011000","00000011",
     "00000001","00001000","01000000","00000011",
     "00000001","00101001","01001000","00000011",
     "00000010","01110011","10011000","00000011",
     "00000011","00011000","11000000","00000011",
     "00000011","00111001","11001000","00000011",
     "00000011","01011010","11010000","00000011",
     "00000011","01111011","11011000","00000011",
     "00011100","00000011","00000000","00111000",
     "00011100","00000100","00000000","00111000",
     "00010100","01100011","00000000","00001000",
     "00000000","01100100","00011000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000100","00011000","00000000","00010000",
     "00011100","00011001","00000000","00111100",
     "00011100","00001000","00000000","00111101",
     "00010101","00001000","00000000","00010000",
     "00000001","00011001","11001000","00000111",
     "00011100","00011010","00000000","00111110",
     "00011100","00001000","00000000","00111111",
     "00010101","00001000","00000000","00010000",
     "00000001","00011010","11010000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000001","00001000","01000000","00000011",
     "00000100","00000100","00000000","00110100",
     "00000001","00101001","01001000","00000011",
     "00000011","10011100","11100000","00000011",
     "00000000","00011001","11100000","00000001",
     "00000100","00010011","00000000","00010000",
     "00101000","00010011","00000000","00000111",
     "00010101","00101001","00000000","00000001",
     "00100111","10000000","00000000","00000011",
     "00010111","10011100","00000000","00000001",
     "00001010","01110011","00000000","00000001",
     "00110000","00000000","00000000","00011101",
     "00010001","00101001","00000000","00000001",
     "00110000","00000000","00000000","00100000",
     "00000011","10011100","11100000","00000011",
     "00000011","10001001","11100000","00000111",
     "00100001","00011100","00000000","00000000",
     "00000101","00001000","00000000","00000001",
     "00100001","00011001","00000000","00000000",
     "00000011","00111010","11001000","00000001",
     "00000101","00001000","00000000","00000001",
     "00100101","00000100","11111111","11101100",
     "00000000","10000100","00100000","00000011",
     "00000001","00001000","01000000","00000011",
     "00000001","00101001","01001000","00000011",
     "00000010","01010010","10010000","00000011",
     "00000010","01110011","10011000","00000011",
     "00000010","10010100","10100000","00000011",
     "00000010","10110101","10101000","00000011",
     "00000010","11010110","10110000","00000011",
     "00000010","11110111","10111000","00000011",
     "00000011","00011000","11000000","00000011",
     "00000011","00111001","11001000","00000011",
     "00000011","01011010","11010000","00000011",
     "00000011","01111011","11011000","00000011",
     "00000011","10011100","11100000","00000011",
     "00000011","10111101","11101000","00000011",
     "00000011","11011110","11110000","00000011",
     "00000011","11111111","11111000","00000011",
     "00000100","00011000","00000000","00011010",
     "00000111","00011000","00000000","00011010",
     "00000111","00011000","00000000","00011010",
     "00000100","00000100","00000000","00000111",
     "00010100","10000100","00000000","00011101",
     "00101011","00000000","00000000","10000001",
     "00001011","00011000","00000000","00000001",
     "00011111","00111101","00000000","00000000",
     "00000000","01111101","11101000","00000101",
     "00010111","10111101","00000000","00010000",
     "00000111","00111001","00000000","00000001",
     "00011111","00101000","00000000","00000000",
     "00001011","00111001","00000000","00000001",
     "00000001","00000011","01000000","00000101",
     "00000001","00011101","11101000","00000111",
     "00000011","10111110","11101000","00000001",
     "00000011","10111111","11101000","00000001",
     "00000000","10011101","01001000","00000101",
     "00010111","10111101","00000000","00000011",
     "00000001","00001000","01000000","00000011",
     "00000010","11110111","10111000","00000011",
     "00000100","00001000","00000000","00100000",
     "00001001","00001000","00000000","00011101",
     "00101001","00000000","00000000","00000111",
     "00010110","11110111","00000000","00000001",
     "00100101","00100000","00000000","00000011",
     "00010101","00101001","00000000","00000001",
     "00001001","00001000","00000000","00000001",
     "00110000","00000000","00000000","01010101",
     "00010010","11110111","00000000","00000001",
     "00110000","00000000","00000000","01011000",
     "00000001","00101001","01001000","00000011",
     "00000001","00110111","01001000","00000111",
     "00000001","00111101","11101000","00000111",
     "00000000","00011101","11110000","00000001",
     "00000010","01010010","10010000","00000011",
     "00000010","01110011","10011000","00000011",
     "00000010","10010100","10100000","00000011",
     "00000000","00011101","10010000","00000001",
     "00000110","01110011","00000000","00010000",
     "00101010","01100000","00000000","00000111",
     "00010110","10010100","00000000","00000001",
     "00100110","01000000","00000000","00000011",
     "00010110","01010010","00000000","00000001",
     "00001010","01110011","00000000","00000001",
     "00110000","00000000","00000000","01100110",
     "00010010","10010100","00000000","00000001",
     "00110000","00000000","00000000","01101001",
     "00000010","01010010","10010000","00000011",
     "00000010","01010100","10010000","00000111",
     "00100011","00110010","00000000","00000000",
     "00000111","00111001","00000000","00000001",
     "00100011","00111101","00000000","00000000",
     "00001011","00111001","00000000","00000001",
     "00000001","00101001","01001000","00000011",
     "00000010","01010010","10010000","00000011",
     "00000010","01110011","10011000","00000011",
     "00000010","10010100","10100000","00000011",
     "00000010","10110101","10101000","00000011",
     "00000010","11010110","10110000","00000011",
     "00000010","11110111","10111000","00000011",
     "00000011","11011111","10010000","00000001",
     "00001110","01010011","00000000","00011111",
     "00000000","00010011","01001000","00000001",
     "00101010","01100000","00000000","00000100",
     "00010110","10110101","00000000","00000001",
     "00010010","10110101","00000000","00000001",
     "00001010","01110011","00000000","00000001",
     "00110000","00000000","00000000","01111110",
     "00000100","00010011","00000000","00100000",
     "00000010","01101001","10011000","00000011",
     "00101010","01100000","00000000","00000011",
     "00010110","10110101","00000000","00000001",
     "00001010","01110011","00000000","00000001",
     "00110000","00000000","00000000","10000101",
     "00011111","01110110","00000000","01000000",
     "00000111","01111011","00000000","00000001",
     "00011111","01110111","00000000","01000000",
     "00000000","01110111","10111000","00000101",
     "00001011","01111011","00000000","00000001",
     "00010110","11010110","00000000","00010000",
     "00000010","11010111","10110000","00000111",
     "00000010","11011110","10110000","00000001",
     "00000010","11011111","10110000","00000001",
     "00000010","01010010","10010000","00000011",
     "00000010","10110110","10010000","00000101",
     "00000001","00001000","01000000","00000011",
     "00000010","10110101","10101000","00000011",
     "00000001","00001001","01000000","00000001",
     "00101001","00000000","00000000","00000111",
     "00010110","10110101","00000000","00000001",
     "00100110","01000000","00000000","00000011",
     "00010110","01010010","00000000","00000001",
     "00001001","00001000","00000000","00000001",
     "00110000","00000000","00000000","10010111",
     "00010010","10110101","00000000","00000001",
     "00110000","00000000","00000000","10011010",
     "00000010","01010010","10010000","00000011",
     "00000010","01010101","10010000","00000111",
     "00101000","00001001","00000000","00000011",
     "00010110","11010110","00000000","00000001",
     "00001001","00101001","00000000","00000001",
     "00110000","00000000","00000000","10100001",
     "00000010","01010110","10110000","00000111",
     "00000000","00010110","11111000","00000001",
     "00000000","00010110","10100000","00000001",
     "00000010","01010010","10010000","00000011",
     "00000010","01110011","10011000","00000011",
     "00000010","10110101","10101000","00000011",
     "00000110","01110011","00000000","00010000",
     "00101010","01100000","00000000","00000111",
     "00010110","10110101","00000000","00000001",
     "00100110","10000000","00000000","00000011",
     "00010110","10010100","00000000","00000001",
     "00001010","01110011","00000000","00000001",
     "00110000","00000000","00000000","10101100",
     "00010010","10110101","00000000","00000001",
     "00110000","00000000","00000000","10101111",
     "00000010","10010100","10100000","00000011",
     "00000010","10010101","10100000","00000111",
     "00100011","01110100","00000000","01000000",
     "00000111","01111011","00000000","00000001",
     "00100011","01110110","00000000","01000000",
     "00001011","01111011","00000000","00000001",
     "00000111","00111001","00000000","00000010",
     "00000011","01011010","11010000","00000011",
     "00001011","00111010","00000000","00110100",
     "00100111","01000000","00000000","00000001",
     "00000011","00111001","11001000","00000011",
     "00000111","01111011","00000000","00000010",
     "00000011","10011100","11100000","00000011",
     "00001011","01111100","00000000","00001000",
     "00100111","10000000","00000000","00000001",
     "00000011","01111011","11011000","00000011",
     "00110000","00000000","00000000","01000011",
     "11111100","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000011",
     "00000000","00100001","00001000","00000011",
     "00000000","01000010","00010000","00000011",
     "00000000","01100011","00011000","00000011",
     "00000000","10000100","00100000","00000011",
     "00011100","00000011","00000000","00111000",
     "00011100","00000100","00000000","00111000",
     "00010100","01100011","00000000","00001000",
     "00000000","01100100","00011000","00000111",
     "00000000","10000100","00100000","00000011",
     "00011100","00000001","00000000","00110100",
     "00010100","00100001","00000000","00010000",
     "00011100","10000100","00000000","00110101",
     "00000000","10000011","00100000","00000101",
     "00000000","00100100","00001000","00000111",
     "00000000","10000100","00100000","00000011",
     "00011100","00000010","00000000","00110110",
     "00010100","01000010","00000000","00010000",
     "00011100","10000100","00000000","00110111",
     "00000000","10000011","00100000","00000101",
     "00000000","01000100","00010000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","10100101","00101000","00000011",
     "00000100","10100101","00000000","00000100",
     "00011100","00000110","00000000","00000000",
     "00010100","11000110","00000000","00010000",
     "00011100","00000100","00000000","00000001",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","00100110","00001000","00000001",
     "00011100","00000110","00000000","00000010",
     "00010100","11000110","00000000","00010000",
     "00011100","00000100","00000000","00000011",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","01000110","00010000","00000001",
     "00000000","00000000","00000000","00000011",
     "00000000","11100111","00111000","00000011",
     "00000100","11100111","00000000","00001100",
     "00000010","00010000","10000000","00000011",
     "00000010","00110001","10001000","00000011",
     "00000000","00100010","10000000","00000101",
     "00000000","00100010","10001000","00001001",
     "00000010","00010001","00001000","00001001",
     "00000001","01101011","01011000","00000011",
     "00000001","01100010","01011000","00000111",
     "00000001","10001100","01100000","00000011",
     "00000001","10000001","01100000","00000111",
     "00000001","11001110","01110000","00000011",
     "00000001","11001011","01110000","00000111",
     "00000001","11101111","01111000","00000011",
     "00000001","11101100","01111000","00000111",
     "00001101","01101011","00000000","00011111",
     "00001101","11001110","00000000","00011111",
     "00101000","00001110","00000000","00000011",
     "00010101","11101111","00000000","00000001",
     "00001001","11001110","00000000","00000001",
     "00101101","11000000","11111111","11111101",
     "00000001","01001010","01010000","00000011",
     "00101001","01100000","00000000","00000111",
     "00010101","01001010","00000000","00000001",
     "00100101","10000000","00000000","00000011",
     "00010101","10001100","00000000","00000001",
     "00001001","01101011","00000000","00000001",
     "00110000","00000000","00000001","00000011",
     "00010001","01001010","00000000","00000001",
     "00110000","00000000","00000001","00000110",
     "00000001","10001100","01100000","00000011",
     "00000001","10001010","01100000","00000111",
     "00000001","10001111","01100000","00000111",
     "00000000","00100001","00001000","00000011",
     "00000000","00101100","00001000","00000111",
     "00011100","10100110","00000000","00000000",
     "00010100","11000110","00000000","00010000",
     "00000100","10100101","00000000","00000001",
     "00011100","10100100","00000000","00000000",
     "00000100","10100101","00000000","00000001",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","00100110","00001000","00000001",
     "00000010","00010000","10000000","00000011",
     "00000010","00110001","10001000","00000011",
     "00000000","00100010","10000000","00000101",
     "00000000","00100010","10001000","00001001",
     "00000010","00010001","00010000","00001001",
     "00000001","01101011","01011000","00000011",
     "00000001","01100001","01011000","00000111",
     "00000001","10001100","01100000","00000011",
     "00000001","10000010","01100000","00000111",
     "00000001","11001110","01110000","00000011",
     "00000001","11001011","01110000","00000111",
     "00000001","11101111","01111000","00000011",
     "00000001","11101100","01111000","00000111",
     "00001101","01101011","00000000","00011111",
     "00001101","11001110","00000000","00011111",
     "00101000","00001110","00000000","00000011",
     "00010101","11101111","00000000","00000001",
     "00001001","11001110","00000000","00000001",
     "00101101","11000000","11111111","11111101",
     "00000001","01001010","01010000","00000011",
     "00101001","01100000","00000000","00000111",
     "00010101","01001010","00000000","00000001",
     "00100101","10000000","00000000","00000011",
     "00010101","10001100","00000000","00000001",
     "00001001","01101011","00000000","00000001",
     "00110000","00000000","00000001","00101101",
     "00010001","01001010","00000000","00000001",
     "00110000","00000000","00000001","00110000",
     "00000001","10001100","01100000","00000011",
     "00000001","10001010","01100000","00000111",
     "00000001","10001111","01100000","00000111",
     "00000000","01000010","00010000","00000011",
     "00000000","01001100","00010000","00000111",
     "00011100","10100110","00000000","00000000",
     "00010100","11000110","00000000","00010000",
     "00000100","10100101","00000000","00000001",
     "00011100","10100100","00000000","00000000",
     "00000100","10100101","00000000","00000001",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","01000110","00010000","00000001",
     "00001000","11100111","00000000","00000001",
     "00101100","00000111","11111111","10101010",
     "11111100","00000000","00000000","00000000",
     "00000000","00000000","00000000","00000011",
     "00000000","00100001","00001000","00000011",
     "00000000","01000010","00010000","00000011",
     "00000000","01100011","00011000","00000011",
     "00000000","10000100","00100000","00000011",
     "00000000","10000100","00100000","00000011",
     "00011100","00000011","00000000","00111000",
     "00011100","00000100","00000000","00111000",
     "00010100","01100011","00000000","00001000",
     "00000000","01100100","00011000","00000111",
     "00000000","10000100","00100000","00000011",
     "00011100","00000001","00000000","00110100",
     "00010100","00100001","00000000","00010000",
     "00011100","10000100","00000000","00110101",
     "00000000","10000011","00100000","00000101",
     "00000000","00100100","00001000","00000111",
     "00000000","10000100","00100000","00000011",
     "00011100","00000010","00000000","00110110",
     "00010100","01000010","00000000","00010000",
     "00011100","10000100","00000000","00110111",
     "00000000","10000011","00100000","00000101",
     "00000000","01000100","00010000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","10100101","00101000","00000011",
     "00000100","10100101","00000000","00110011",
     "00000000","00000000","00000000","00000011",
     "00000000","11100111","00111000","00000011",
     "00000100","11100111","00000000","00001100",
     "00011100","10100110","00000000","00000000",
     "00000000","11000011","00110000","00000101",
     "00001000","10100101","00000000","00000001",
     "00011100","10100100","00000000","00000000",
     "00010100","10000100","00000000","00010000",
     "00001000","10100101","00000000","00000001",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","01000110","00010000","00000011",
     "00000010","01010010","10010000","00000011",
     "00000010","01110011","10011000","00000011",
     "00000000","00110011","10011000","00000111",
     "00000000","01010010","10010000","00000111",
     "00001110","01110011","00000000","00011111",
     "00000000","00000000","00000000","00000011",
     "00000010","10010100","10100000","00000011",
     "00000010","10110101","10101000","00000011",
     "00000010","11010110","10110000","00000011",
     "00000010","11110111","10111000","00000011",
     "00101000","00010011","00000000","00010111",
     "00000000","00010011","10100000","00000001",
     "00010110","10110101","00000000","00000001",
     "00010010","10110101","00000000","00000001",
     "00001010","10010100","00000000","00000001",
     "00101100","00010100","11111111","11111100",
     "00000010","01010101","10101000","00000101",
     "00000010","01110100","10100000","00000001",
     "00000110","11110111","00000000","00100000",
     "00000010","11110011","10011000","00000011",
     "00101000","00010011","00000000","00000111",
     "00010110","11010110","00000000","00000001",
     "00100110","01000000","00000000","00000011",
     "00010110","01010010","00000000","00000001",
     "00001010","01110011","00000000","00000001",
     "00110000","00000000","00000001","01111111",
     "00010010","11010110","00000000","00000001",
     "00110000","00000000","00000001","10000010",
     "00000010","01010010","10010000","00000011",
     "00000010","11110100","10100000","00000011",
     "00010110","10110101","00000000","00000001",
     "00001010","10010100","00000000","00000001",
     "00101100","00010100","11111111","11111101",
     "00000010","10110110","10010000","00000111",
     "00000000","01000010","00010000","00000011",
     "00000000","01010010","00010000","00000111",
     "00000010","00010000","10000000","00000011",
     "00000010","00110001","10001000","00000011",
     "00000000","00100010","10000000","00000101",
     "00000000","00100010","10001000","00001001",
     "00000010","00010001","00010000","00001001",
     "00011100","10100110","00000000","00000000",
     "00000000","11000011","00110000","00000101",
     "00001000","10100101","00000000","00000001",
     "00011100","10100100","00000000","00000000",
     "00010100","10000100","00000000","00010000",
     "00001000","10100101","00000000","00000001",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","00100110","00001000","00000011",
     "00000010","01010010","10010000","00000011",
     "00000010","01110011","10011000","00000011",
     "00000000","00110010","10010000","00000111",
     "00000000","01010011","10011000","00000111",
     "00001110","01110011","00000000","00011111",
     "00000000","00000000","00000000","00000011",
     "00000010","10010100","10100000","00000011",
     "00000010","10110101","10101000","00000011",
     "00000010","11010110","10110000","00000011",
     "00000010","11110111","10111000","00000011",
     "00101000","00010011","00000000","00010111",
     "00000000","00010011","10100000","00000001",
     "00010110","10110101","00000000","00000001",
     "00010010","10110101","00000000","00000001",
     "00001010","10010100","00000000","00000001",
     "00101100","00010100","11111111","11111100",
     "00000010","01010101","10101000","00000101",
     "00000010","01110100","10100000","00000001",
     "00000110","11110111","00000000","00100000",
     "00000010","11110011","10011000","00000011",
     "00101000","00010011","00000000","00000111",
     "00010110","11010110","00000000","00000001",
     "00100110","01000000","00000000","00000011",
     "00010110","01010010","00000000","00000001",
     "00001010","01110011","00000000","00000001",
     "00110000","00000000","00000001","10110001",
     "00010010","11010110","00000000","00000001",
     "00110000","00000000","00000001","10110100",
     "00000010","01010010","10010000","00000011",
     "00000010","11110100","10100000","00000011",
     "00010110","10110101","00000000","00000001",
     "00001010","10010100","00000000","00000001",
     "00101100","00010100","11111111","11111101",
     "00000010","10110110","10010000","00000111",
     "00000000","00100001","00001000","00000011",
     "00000000","00110010","00001000","00000111",
     "00000010","00010000","10000000","00000011",
     "00000010","00110001","10001000","00000011",
     "00000000","00100010","10000000","00000101",
     "00000000","00100010","10001000","00001001",
     "00000010","00010001","00001000","00001001",
     "00001000","11100111","00000000","00000001",
     "00101100","00000111","11111111","10011010",
     "00000000","10000100","00100000","00000011",
     "00011100","00000110","00000000","00000000",
     "00010100","11000110","00000000","00010000",
     "00011100","00000100","00000000","00000001",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","00100110","00001000","00000011",
     "00011100","00000110","00000000","00000010",
     "00010100","11000110","00000000","00010000",
     "00011100","00000100","00000000","00000011",
     "00000000","10000011","00100000","00000101",
     "00000000","11000100","00110000","00000111",
     "00000000","10000100","00100000","00000011",
     "00000000","01000110","00010000","00000011",
     "11111100","00000000","00000000","00000000"
      );  
    begin
        out_imem <= rom_data(to_integer(unsigned(in_pc(31 downto 0)))) & rom_data(to_integer(unsigned(in_pc(31 downto 0)) + 1 )) & rom_data(to_integer(unsigned(in_pc(31 downto 0)) + 2 )) & rom_data(to_integer(unsigned(in_pc(31 downto 0)) + 3 ));
end Behavioral;

